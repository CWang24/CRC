`timescale 1ns/10ps
module tb;
reg [7:0] data_in;
crc crc_tb(data_in,crc_out);
initial
	begin
	data_in=8'b11111111;
	#2;
	data_in=8'b00000000;
	#2;
	data_in=8'b00000001;
	#2;
	data_in=8'b00000010;
	#2;
	data_in=8'b00000011;
	#2;
	data_in=8'b00000100;
	#2;
	data_in=8'b00000101;
	#2;
	data_in=8'b00000110;
	#2;
	data_in=8'b00000111;
	#2;
	data_in=8'b00001000;
	#2;
	data_in=8'b00001001;
	#2;
	data_in=8'b00001010;
	#2;
	data_in=8'b00001011;
	#2;
	data_in=8'b00001100;
	#2;
	data_in=8'b00001101;
	#2;
	data_in=8'b00001110;
	#2;
	data_in=8'b00001111;
	#2;
	data_in=8'b00010000;
	#2;
	data_in=8'b00010001;
	#2;
	data_in=8'b00010010;
	#2;
	data_in=8'b00010011;
	#2;
	data_in=8'b00010100;
	#2;
	data_in=8'b00010101;
	#2;
	data_in=8'b00010110;
	#2;
	data_in=8'b00010111;
	#2;
	data_in=8'b00011000;
	#2;
	data_in=8'b00011001;
	#2;
	data_in=8'b00011010;
	#2;
	data_in=8'b00011011;
	#2;
	data_in=8'b00011100;
	#2;
	data_in=8'b00011101;
	#2;
	data_in=8'b00011110;
	#2;
	data_in=8'b00011111;
	#2;
	data_in=8'b00100000;
	#2;
	data_in=8'b00100001;
	#2;
	data_in=8'b00100010;
	#2;
	data_in=8'b00100011;
	#2;
	data_in=8'b00100100;
	#2;
	data_in=8'b00100101;
	#2;
	data_in=8'b00100110;
	#2;
	data_in=8'b00100111;
	#2;
	data_in=8'b00101000;
	#2;
	data_in=8'b00101001;
	#2;
	data_in=8'b00101010;
	#2;
	data_in=8'b00101011;
	#2;
	data_in=8'b00101100;
	#2;
	data_in=8'b00101101;
	#2;
	data_in=8'b00101110;
	#2;
	data_in=8'b00101111;
	#2;
	data_in=8'b00110000;
	#2;
	data_in=8'b00110001;
	#2;
	data_in=8'b00110010;
	#2;
	data_in=8'b00110011;
	#2;
	data_in=8'b00110100;
	#2;
	data_in=8'b00110101;
	#2;
	data_in=8'b00110110;
	#2;
	data_in=8'b00110111;
	#2;
	data_in=8'b00111000;
	#2;
	data_in=8'b00111001;
	#2;
	data_in=8'b00111010;
	#2;
	data_in=8'b00111011;
	#2;
	data_in=8'b00111100;
	#2;
	data_in=8'b00111101;
	#2;
	data_in=8'b00111110;
	#2;
	data_in=8'b00111111;
	#2;
	data_in=8'b01000000;
	#2;
	data_in=8'b01000001;
	#2;
	data_in=8'b01000010;
	#2;
	data_in=8'b01000011;
	#2;
	data_in=8'b01000100;
	#2;
	data_in=8'b01000101;
	#2;
	data_in=8'b01000110;
	#2;
	data_in=8'b01000111;
	#2;
	data_in=8'b01001000;
	#2;
	data_in=8'b01001001;
	#2;
	data_in=8'b01001010;
	#2;
	data_in=8'b01001011;
	#2;
	data_in=8'b01001100;
	#2;
	data_in=8'b01001101;
	#2;
	data_in=8'b01001110;
	#2;
	data_in=8'b01001111;
	#2;
	data_in=8'b01010000;
	#2;
	data_in=8'b01010001;
	#2;
	data_in=8'b01010010;
	#2;
	data_in=8'b01010011;
	#2;
	data_in=8'b01010100;
	#2;
	data_in=8'b01010101;
	#2;
	data_in=8'b01010110;
	#2;
	data_in=8'b01010111;
	#2;
	data_in=8'b01011000;
	#2;
	data_in=8'b01011001;
	#2;
	data_in=8'b01011010;
	#2;
	data_in=8'b01011011;
	#2;
	data_in=8'b01011100;
	#2;
	data_in=8'b01011101;
	#2;
	data_in=8'b01011110;
	#2;
	data_in=8'b01011111;
	#2;
	data_in=8'b01100000;
	#2;
	data_in=8'b01100001;
	#2;
	data_in=8'b01100010;
	#2;
	data_in=8'b01100011;
	#2;
	data_in=8'b01100100;
	#2;
	data_in=8'b01100101;
	#2;
	data_in=8'b01100110;
	#2;
	data_in=8'b01100111;
	#2;
	data_in=8'b01101000;
	#2;
	data_in=8'b01101001;
	#2;
	data_in=8'b01101010;
	#2;
	data_in=8'b01101011;
	#2;
	data_in=8'b01101100;
	#2;
	data_in=8'b01101101;
	#2;
	data_in=8'b01101110;
	#2;
	data_in=8'b01101111;
	#2;
	data_in=8'b01110000;
	#2;
	data_in=8'b01110001;
	#2;
	data_in=8'b01110010;
	#2;
	data_in=8'b01110011;
	#2;
	data_in=8'b01110100;
	#2;
	data_in=8'b01110101;
	#2;
	data_in=8'b01110110;
	#2;
	data_in=8'b01110111;
	#2;
	data_in=8'b01111000;
	#2;
	data_in=8'b01111001;
	#2;
	data_in=8'b01111010;
	#2;
	data_in=8'b01111011;
	#2;
	data_in=8'b01111100;
	#2;
	data_in=8'b01111101;
	#2;
	data_in=8'b01111110;
	#2;
	data_in=8'b01111111;
	#2;
	data_in=8'b10000000;
	#2;
	data_in=8'b10000001;
	#2;
	data_in=8'b10000010;
	#2;
	data_in=8'b10000011;
	#2;
	data_in=8'b10000100;
	#2;
	data_in=8'b10000101;
	#2;
	data_in=8'b10000110;
	#2;
	data_in=8'b10000111;
	#2;
	data_in=8'b10001000;
	#2;
	data_in=8'b10001001;
	#2;
	data_in=8'b10001010;
	#2;
	data_in=8'b10001011;
	#2;
	data_in=8'b10001100;
	#2;
	data_in=8'b10001101;
	#2;
	data_in=8'b10001110;
	#2;
	data_in=8'b10001111;
	#2;
	data_in=8'b10010000;
	#2;
	data_in=8'b10010001;
	#2;
	data_in=8'b10010010;
	#2;
	data_in=8'b10010011;
	#2;
	data_in=8'b10010100;
	#2;
	data_in=8'b10010101;
	#2;
	data_in=8'b10010110;
	#2;
	data_in=8'b10010111;
	#2;
	data_in=8'b10011000;
	#2;
	data_in=8'b10011001;
	#2;
	data_in=8'b10011010;
	#2;
	data_in=8'b10011011;
	#2;
	data_in=8'b10011100;
	#2;
	data_in=8'b10011101;
	#2;
	data_in=8'b10011110;
	#2;
	data_in=8'b10011111;
	#2;
	data_in=8'b10100000;
	#2;
	data_in=8'b10100001;
	#2;
	data_in=8'b10100010;
	#2;
	data_in=8'b10100011;
	#2;
	data_in=8'b10100100;
	#2;
	data_in=8'b10100101;
	#2;
	data_in=8'b10100110;
	#2;
	data_in=8'b10100111;
	#2;
	data_in=8'b10101000;
	#2;
	data_in=8'b10101001;
	#2;
	data_in=8'b10101010;
	#2;
	data_in=8'b10101011;
	#2;
	data_in=8'b10101100;
	#2;
	data_in=8'b10101101;
	#2;
	data_in=8'b10101110;
	#2;
	data_in=8'b10101111;
	#2;
	data_in=8'b10110000;
	#2;
	data_in=8'b10110001;
	#2;
	data_in=8'b10110010;
	#2;
	data_in=8'b10110011;
	#2;
	data_in=8'b10110100;
	#2;
	data_in=8'b10110101;
	#2;
	data_in=8'b10110110;
	#2;
	data_in=8'b10110111;
	#2;
	data_in=8'b10111000;
	#2;
	data_in=8'b10111001;
	#2;
	data_in=8'b10111010;
	#2;
	data_in=8'b10111011;
	#2;
	data_in=8'b10111100;
	#2;
	data_in=8'b10111101;
	#2;
	data_in=8'b10111110;
	#2;
	data_in=8'b10111111;
	#2;
	data_in=8'b11000000;
	#2;
	data_in=8'b11000001;
	#2;
	data_in=8'b11000010;
	#2;
	data_in=8'b11000011;
	#2;
	data_in=8'b11000100;
	#2;
	data_in=8'b11000101;
	#2;
	data_in=8'b11000110;
	#2;
	data_in=8'b11000111;
	#2;
	data_in=8'b11001000;
	#2;
	$stop; 
	end
endmodule
